`define DATA_WIDTH 32
`define AL_SIZE 64
`define NUM_CHECKPOINTS 16
`define NUM_BRANCHES_RESOLVED 2
`define ADDR_WIDTH 32
`define NUM_INSTRS_COMPLETED 2
`define INSTR_MEM_SIZE 1024
`define DATA_MEM_SIZE 16
`define NUM_WRITES_CORE 1
`define NUM_ARITH_CORE 2

import riscv_pkg::*;