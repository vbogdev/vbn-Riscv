`define DATA_WIDTH 32
`define ADDR_WIDTH 32
`define INSTR_MEM_SIZE 1024
`define DATA_MEM_SIZE 16
`define NUM_WRITES_CORE 1
`define NUM_CORES 2

import riscv_pkg::*;